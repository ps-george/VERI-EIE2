module starting_line_fsm(



);



endmodule
